Library IEEE;
use IEEE.std_logic_1164.all;


ENTITY TP_Base_addition IS
port( 
A1,B1,Cin : in std_logic;			 
S,Cout:out std_logic
);
END TP_Base_addition;

architecture ar of TP_Base_addition is
BEGIN



END ar ;